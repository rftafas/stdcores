----------------------------------------------------------------------------------------------------------
-- Simple Serial Controllers - SPI MASTER
-- Ricardo Tafas
-- This is open source code licensed under LGPL.
-- By using it on your system you agree with all LGPL conditions.
-- This code is provided AS IS, without any sort of warranty.
-- Author: Ricardo F Tafas Jr
-- 2020
---------------------------------------------------------------------------------------------------------
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;
library expert;
  use expert.std_logic_expert.all;
library stdblocks;
  use stdblocks.sync_lib.all;
library stdcores;
	use stdcores.axis_s_spim_pkg.all;


entity axis_s_spi_m_tb is
end axis_s_spi_m_tb;

architecture simulation of axis_s_spi_m_tb is


begin

end behavioral;
